/****************************************
*****************************************
|------	AStarSim v1.2 ------------------|
|------	By Tristan Michael -------------|
*****************************************
|------	Started: 5/08/04 ---------------|
|------	Updated: 5/25/04 ---------------|
*****************************************
*****************************************/

//---------------------------------------
//---------------------------------------
//GLOBALS
//---------------------------------------

//----A* Algorithm specific Variables

//width and height in tiles +1
#define TIMEOUT 1000
#define MAP_WIDTH 1001
#define MAP_HEIGHT 1001
#define MAX_OPEN 9999
#define H_D 10 //used when calculating H
#define G_D 10 //used when calculating G
#define GC_D 14 //used when calculating G at a corner
#define TILES 1 //number of tiles to use in a node(1 = 1X1 nodes and 16X16 tiles, 2 = 2X2 nodes and 32x32 tiles) 

//defines for determining 'which'
#define NODE_NONE 0
#define NODE_OPEN 1 
#define NODE_CLOSED 2

//individual node properties
int node_which[MAP_WIDTH][MAP_HEIGHT];
int node_G[MAP_WIDTH][MAP_HEIGHT];
int node_H[MAP_WIDTH][MAP_HEIGHT];
int node_cost[MAP_WIDTH][MAP_HEIGHT];
int node_parentX[MAP_WIDTH][MAP_HEIGHT];
int node_parentY[MAP_WIDTH][MAP_HEIGHT];
int nAStartStartTime;

struct plot{
	int x;
	int y;
}

//Active nodes used to keep tract of what nodes to pay attention to.
int activeNodes;
plot activeList[MAX_OPEN];

int open;
int openList[MAX_OPEN];

int paths;
plot path[MAX_OPEN]; //result of findPath();

//------------------------------------------------
//MAIN CODE
//------------------------------------------------
//Finds path using A* algorithm
//0=error
plot temp;
plot cur;
int timeTrack;

int findPath(int ent, int x1, int y1, int x2, int y2){
	int i, chkValue, foundPath, tempIndex, tempCost;
//Check for immediate errors in path
	if(x1 == x2 && y1 == y2){
		log("EXIT: already at target position");
		return 0;
	}
	if(chkObs(x2,y2)){
		log("EXIT: target is an obstruction");
		return 0;
	}
	//timer=0;
	nAStartStartTime = timer;
	
//set-up initial variables
	cur.x=x2;
	cur.y=y2;
	
	paths=0;
	open=0;
	
	activeNodes=1;
	activeList[activeNodes].x=cur.x;
	activeList[activeNodes].y=cur.y;
	
	node_which[cur.x][cur.y]=NODE_OPEN;
	node_G[cur.x][cur.y]=0;
	node_H[cur.x][cur.y]=H_D*(abs(cur.x-x1) + abs(cur.y-y1));
	node_Cost[cur.x][cur.y]=node_G[cur.x][cur.y] + node_H[cur.x][cur.y];
	node_parentX[cur.x][cur.y]=x2;
	node_parentY[cur.x][cur.y]=y2;
	
	addOpenID(activeNodes);

//----Start Loop
	while(!foundPath){		
		if(open == 0){
			log("EXIT: Couldent find another open node, no path.");
			return(0); //No path
		}
		if(timer > TIMEOUT+nAStartStartTime){
			log("EXIT: Timeout.");
			return(0);
		}
//#2. add lowest open to closed list and set as current

	//DEBUG
		line(activeList[openList[1]].x*(16*TILES)+8-xwin, activeList[openList[1]].y*(16*TILES)+8-ywin, node_parentX[activeList[openList[1]].x][activeList[openList[1]].y]*(16*TILES)+8-xwin, node_parentY[activeList[openList[1]].x][activeList[openList[1]].y]*(16*TILES)+8-ywin, RGB(0,0,255), screen);
		rect(activeList[openList[1]].x*(16*TILES)-xwin, activeList[openList[1]].y*(16*TILES)-ywin, activeList[openList[1]].x*(16*TILES)+(16*TILES)-xwin, activeList[openList[1]].y*(16*TILES)+(16*TILES)-ywin, RGB(255,0,0), screen);		
	//DEBUG
		
		cur.x=activeList[openList[1]].x;
		cur.y=activeList[openList[1]].y;
		node_which[cur.x][cur.y]=NODE_CLOSED;
		
		closeOpenID(1);

//#3. find adjacent squares and add to open list
		for(temp.y=cur.y-1;temp.y<=cur.y+1;temp.y++)
		if( !chkObs(cur.x,temp.y) ) //diagonal correction (top/bottom)
		for(temp.x=cur.x-1;temp.x<=cur.x+1;temp.x++)
		if( !chkObs(temp.x, temp.y-(temp.y-cur.y)) ) //diagonal correction
		if(!chkObs(temp.x, temp.y)){
		
		//look up node type
			chkValue=activeChk(temp.x, temp.y);
			
		//figure out path movement cost
			if(abs(temp.x-cur.x) == 1 && abs(temp.y-cur.y) == 1) tempCost=GC_D;
			else tempCost=G_D;
			
		//add new nodes
			if(chkValue == NODE_NONE){
				if(activeNodes == MAX_OPEN-1){
					log("EXIT: path too long");
					return(0);
				}
				activeNodes++;
				activeList[activeNodes].x=temp.x;
				activeList[activeNodes].y=temp.y;

				node_which[temp.x][temp.y]=NODE_OPEN;
				
				node_G[temp.x][temp.y]=node_G[cur.x][cur.y]+tempCost;
				node_H[temp.x][temp.y]=H_D*(abs(temp.x-x1) + abs(temp.y-y1));
				node_cost[temp.x][temp.y]=node_G[temp.x][temp.y] + node_H[temp.x][temp.y];
				node_parentX[temp.x][temp.y]=cur.x;
				node_parentY[temp.x][temp.y]=cur.y;	

				addOpenID(activeNodes);
			//DEBUG
				line(temp.x*(16*TILES)+8, temp.y*(16*TILES)+8, cur.x*(16*TILES)+8, cur.y*(16*TILES)+8, RGB(0,0,255), screen);
				rect(temp.x*(16*TILES)-xwin,temp.y*(16*TILES)-ywin,temp.x*(16*TILES)+(16*TILES)-xwin,temp.y*(16*TILES)+(16*TILES)-ywin, RGB(0,255,0), screen);
				printstring(temp.x*(16*TILES)-xwin,temp.y*(16*TILES)-ywin,screen, 0, str(node_cost[temp.x][temp.y]));
				showpage();
			//DEBUG
			}
		//Check already open adjacent nodes to see if current path is better
			else if(chkValue == NODE_OPEN && node_G[temp.x][temp.y] > node_G[cur.x][cur.y]+tempCost){
				node_G[temp.x][temp.y]=node_G[cur.x][cur.y]+tempCost;
				node_cost[temp.x][temp.y]=node_G[temp.x][temp.y] + node_H[temp.x][temp.y];
				node_parentX[temp.x][temp.y]=cur.x;
				node_parentY[temp.x][temp.y]=cur.y;
				
				//line(temp.x*(16*TILES)+8-xwin, temp.y*(16*TILES)+8-ywin, cur.x*(16*TILES)+8-xwin, cur.y*(16*TILES)+8-ywin, RGB(255,0,255), screen);

				chkOpenID( openListChk(temp.x,temp.y) );
			}
		//FOUND TARGET! w00t!!
			if(temp.x == x1 && temp.y == y1){
				foundPath=1;
				cur.x=activeList[openList[1]].x;
				cur.y=activeList[openList[1]].y;
			}
	
		}
//-End loop if path has been found-
	}
//#4. Trace path back from target
	while(cur.x != x2 || cur.y != y2 && paths < MAX_OPEN-1){
		//settile(cur.x,cur.y,0,5);
		
		paths++;
		path[paths].x=cur.x;
		path[paths].y=cur.y;
		
		temp.x=cur.x;
		temp.y=cur.y;
		
		cur.x=node_ParentX[temp.x][temp.y];
		cur.y=node_ParentY[temp.x][temp.y]; 
	}
	//settile(cur.x,cur.y,0,5);
	paths++;
	path[paths].x=cur.x;
	path[paths].y=cur.y;

	temp.x=cur.x;
	temp.y=cur.y;

	cur.x=node_ParentX[temp.x][temp.y];
	cur.y=node_ParentY[temp.x][temp.y]; 
	
//-DONE!
	writePath();
	timeTrack=timer;

	entityMove(ent, entPath);
	
	return(1);
}

//---------------------------------------------------------------
//looks into the active array to find if node[x][y] is active
//0=not active
//1=open
//2=closed
int activeChk(int x, int y){
	int i;
	for(i=1;i<=activeNodes;i++){
		if(activeList[i].x == x && activeList[i].y == y){
			return(node_which[x][y]);
		}
	}
	return(0);
}

int openListChk(int x, int y){
	int i;
	for(i=1;i<=open;i++){
		if(activeList[openList[i]].x == x && activeList[openList[i]].y == y){
			return(i);
		}
	}
	return(0);
}


//note: include entities and map restrictions in obstruction chk
int chkObs(int x, int y){
	int tx,ty;
	x=x*TILES;
	y=y*TILES;
	if (temp.x >= 0 && temp.y >= 0 && temp.x != MAP_WIDTH && temp.y != MAP_HEIGHT){
		for(ty=y;ty<=y+TILES-1;ty++)
		for(tx=x;tx<=x+TILES-1;tx++)
			if(getObs(tx,ty)){
				//rect(tx*(16)-xwin,ty*(16)-ywin,tx*(16)-xwin+(16),ty*(16)-ywin+(16),RGB(255,255,255),screen);
				return(1);
			}
			//else rect(tx*(16)-xwin,ty*(16)-ywin,tx*(16)-xwin+(16),ty*(16)-ywin+(16),0,screen);
	}
	else return(1);
	return(0);
}

//-----------------------------------------------------------------
string entPath;
void writePath(){
	int pastPath;
	entPath="";
	
	for(pastPath=1;pastPath<paths;pastPath++){
			if(path[pastPath].x < path[pastpath+1].x) entPath=entpath+"R"+str(TILES); // right
		else 	if(path[pastPath].x > path[pastpath+1].x) entPath=entpath+"L"+str(TILES); // left
			if(path[pastPath].y < path[pastpath+1].y) entPath=entpath+"D"+str(TILES); // down
		else 	if(path[pastPath].y > path[pastpath+1].y) entPath=entpath+"U"+str(TILES); // up
	}
}

/*int processPath(int e){
	if(!entity.movecode[e] && strCmp(entPath,"") != 0){
		entityMove(e, entPath);
		return(1);
	}
	else if(entity.movecode[e] && strCmp(entPath,"") != 0){
		entPath="";	
	}
	return(0);
}*/

//------------------------------------------------------------
//binary-heap opimization code

void addOpenID(int actIndex){
	int tempOpen;
	open++;
	openList[open]=actIndex;
	int lvl=open;
	
	while(lvl > 1){
		if( node_cost[ activeList[openList[ lvl ]].x ][ activeList[openList[ lvl ]].y ] <= node_cost[ activeList[openList[ lvl/2 ]].x ][ activeList[openList[ lvl/2 ]].y ] ){			tempOpen=openList[lvl/2];
			openList[lvl/2]=openList[lvl];
			openList[lvl]=tempOpen;
			lvl=lvl/2;
		}
		else return;
	}
}

void chkOpenID(int openIndex){
	int tempOpen;
	int lvl=openIndex;
	
	while(lvl > 1){
		if( node_cost[ activeList[openList[ lvl ]].x ][ activeList[openList[ lvl ]].y ] < node_cost[ activeList[openList[ lvl/2 ]].x ][ activeList[openList[ lvl/2 ]].y ] ){			tempOpen=openList[lvl/2];
			openList[lvl/2]=openList[lvl];
			openList[lvl]=tempOpen;
			lvl=lvl/2;
		}
		else return;
	}
}

void closeOpenID(int lvl){
	int tempOpen=openList[open];
	open--;
	openList[1]=tempOpen;
	
	int tempLvl=lvl;
	
	while(1){
	//find lower of the two children
		if( 2*lvl <= open ) //if 1 child exists
			if( node_cost[ activeList[openList[ lvl ]].x ][ activeList[openList[ lvl ]].y ] >= node_cost[ activeList[openList[ lvl*2 ]].x ][ activeList[openList[ lvl*2 ]].y ] )
				tempLvl=lvl*2;
		if(2*lvl+1 <= open) // if both children exist
			if( node_cost[ activeList[openList[ tempLvl ]].x ][ activeList[openList[ tempLvl ]].y ] >= node_cost[ activeList[openList[ lvl*2+1 ]].x ][ activeList[openList[ lvl*2+1 ]].y ] )
				tempLvl=lvl*2+1;
	//swapping
		if(tempLvl != lvl){
			tempOpen=openList[tempLvl];
			openList[tempLvl]=openList[lvl];
			openList[lvl]=tempOpen;
			lvl=tempLvl;
		}
		else return;
	}
}
